`ifdef __EXU_EXU_TOP_V__

module exu_top_module ( 
    input                                               i_csr_trap_flush,
    input   [1                                  : 0]    i_csr_rv_mode,
    input   [`CSR_SATP_WIDTH - 1                : 0]    i_csr_mmu_satp,


    input                                               i_rsv_exu_vld_0,
    input                                               i_rsv_exu_src1_vld_0,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src1_dat_0,
    input                                               i_rsv_exu_src2_vld_0,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src2_dat_0,
    input                                               i_rsv_exu_src3_vld_0,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src3_dat_0,
    input                                               i_rsv_exu_dst_vld_0,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_dst_code_0,
    input   [`IMM_WIDTH - 1                     : 0]    i_rsv_exu_imm_0,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_rsv_exu_rob_id_0,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_rsv_exu_decinfo_bus_0,
    input                                               i_rsv_exu_len_0,
    input   [`CORE_PC_WIDTH - 1                 : 0]    i_rob_exu_addr_0,
    input   [`EXCEPTION_CODE_WIDTH - 1          : 0]    i_rsv_exu_excp_code_0,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_csr_exu_rdat_0,

    input                                               i_rsv_exu_vld_1,
    input                                               i_rsv_exu_src1_vld_1,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src1_dat_1,
    input                                               i_rsv_exu_src2_vld_1,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src2_dat_1,
    input                                               i_rsv_exu_src3_vld_1,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src3_dat_1,
    input                                               i_rsv_exu_dst_vld_1,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_dst_code_1,
    input   [`IMM_WIDTH - 1                     : 0]    i_rsv_exu_imm_1,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_rsv_exu_rob_id_1,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_rsv_exu_decinfo_bus_1,
    input   [`PREDINFO_WIDTH - 1                : 0]    i_rsv_exu_predinfo_bus_1,
    input                                               i_rsv_exu_len_1,
    input   [`CORE_PC_WIDTH - 1                 : 0]    i_rob_exu_addr_1,
    input   [`CORE_PC_WIDTH - 1                 : 0]    i_rob_exu_taddr_1,
    input   [`EXCEPTION_CODE_WIDTH - 1          : 0]    i_rsv_exu_excp_code_1,

    input                                               i_rsv_exu_vld_2,
    input                                               i_rsv_exu_src1_vld_2,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src1_dat_2,
    input                                               i_rsv_exu_src2_vld_2,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src2_dat_2,
    input                                               i_rsv_exu_src3_vld_2,
    input   [`PRF_DATA_WIDTH - 1                : 0]    i_rsv_exu_src3_dat_2,
    input                                               i_rsv_exu_dst_vld_2,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_dst_code_2,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_rsv_exu_decinfo_bus_2,
    input   [`EXCEPTION_CODE_WIDTH - 1          : 0]    i_rsv_exu_excp_code_2,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_rsv_exu_rob_id_2,

    input                                               i_rsv_exu_vld_3,
    input                                               i_rsv_exu_src1_vld_3,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_src1_dat_3,
    input                                               i_rsv_exu_src2_vld_3,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_src2_dat_3,
    input                                               i_rsv_exu_src3_vld_3,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_src3_dat_3,
    input                                               i_rsv_exu_dst_vld_3,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_rsv_exu_dst_code_3,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_rsv_exu_rob_id_3,
    input                                               i_rsv_exu_ld_vld_3,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rsv_exu_ld_id_3,
    input                                               i_rsv_exu_st_vld_3,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_rsv_exu_st_id_3,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_rsv_exu_decinfo_bus_3,
    input   [`IMM_WIDTH - 1                     : 0]    i_rsv_exu_imm_3,
    input   [3                                  : 0]    i_dsp_rsv_vld,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_dsp_rsv_rob_id_0,
    input                                               i_dsp_rsv_ld_vld_0,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_ld_id_0,
    input                                               i_dsp_rsv_st_vld_0,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_st_id_0,
    input                                               i_dsp_rsv_dst_vld_0,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_dsp_rsv_dst_code_0,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_dsp_rsv_decinfo_bus_0,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_dsp_rsv_rob_id_1,
    input                                               i_dsp_rsv_ld_vld_1,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_ld_id_1,
    input                                               i_dsp_rsv_st_vld_1,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_st_id_1,
    input                                               i_dsp_rsv_dst_vld_1,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_dsp_rsv_dst_code_1,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_dsp_rsv_decinfo_bus_1,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_dsp_rsv_rob_id_2,
    input                                               i_dsp_rsv_ld_vld_2,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_ld_id_2,
    input                                               i_dsp_rsv_st_vld_2,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_st_id_2,
    input                                               i_dsp_rsv_dst_vld_2,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_dsp_rsv_dst_code_2,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_dsp_rsv_decinfo_bus_2,
    input   [`ROB_ID_WIDTH - 1                  : 0]    i_dsp_rsv_rob_id_3,
    input                                               i_dsp_rsv_ld_vld_3,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_ld_id_3,
    input                                               i_dsp_rsv_st_vld_3,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_dsp_rsv_st_id_3,
    input                                               i_dsp_rsv_dst_vld_3,
    input   [`PRF_CODE_WIDTH - 1                : 0]    i_dsp_rsv_dst_code_3,
    input   [`DECINFO_WIDTH - 1                 : 0]    i_dsp_rsv_decinfo_bus_3,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_dsp_exu_ld_dsp_ptr,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_dsp_exu_ld_ret_ptr,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_dsp_exu_st_dsp_ptr,
    input   [`SBUFF_ID_WIDTH - 1                : 0]    i_dsp_exu_st_ret_ptr,
    input   [`SBUfF_ID_WIDTH - 1                : 0]    i_dsp_exu_st_ret_cptr,
    input   [3                                  : 0]    i_rob_exu_ret_vld,
    input                                               i_rob_exu_ret_ld_vld_0,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_ld_id_0,
    input                                               i_rob_exu_ret_st_vld_0,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_st_id_0,
    input                                               i_rob_exu_ret_ld_vld_1,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_ld_id_1,
    input                                               i_rob_exu_ret_st_vld_1,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_st_id_1,
    input                                               i_rob_exu_ret_ld_vld_2,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_ld_id_2,
    input                                               i_rob_exu_ret_st_vld_2,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_st_id_2,
    input                                               i_rob_exu_ret_ld_vld_3,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_ld_id_3,
    input                                               i_rob_exu_ret_st_vld_3,
    input   [`LBUFF_ID_WIDTH - 1                : 0]    i_rob_exu_ret_st_id_3,
    input   [`CORE_PC_WIDTH - 1                 : 0]    i_rob_exu_ls_addr,
    input                                               i_rob_dtlb_flush,
    input   [31                                 : 0]    i_rob_dtlb_src1,
    input   [31                                 : 0]    i_rob_dtlb_src2,
    input                                               i_mmu_busy,
    input                                               i_mmu_dtlb_vld,
    input   [`DTLB_TLB_WIDTH - 1                : 0]    i_mmu_dtlb_tlb,
    input   [2                                  : 0]    i_mmu_dtlb_excp_code,
    input                                               i_mmu_dcache_vld,
    input   [`DCACHE_DATA_WIDTH - 1             : 0]    i_mmu_dcache_dat,
    input                                               i_mmu_exu_done,

    output  [`CSR_ADDR_WIDTH - 1                : 0]    o_exu_csr_addr,
    output                                              o_exu_csr_wren,
    output  [`PRF_DATA_WIDTH - 1                : 0]    o_exu_csr_wdat,

    output                                              o_exu_rsv_wren_0,
    output  [`PRF_CODE_WIDTH - 1                : 0]    o_exu_rsv_wr_prf_code_0,
    output  [`PRF_DATA_WIDTH - 1                : 0]    o_exu_rsv_wr_dat_0,
    output                                              o_exu_rsv_busy_0,
    output                                              o_exu_rob_vld_0,
    output  [`EXCEPTION_CODE_WIDTH - 1          : 0]    o_exu_rob_excp_code_0,
    output                                              o_exu_rob_done_0,
    output  [`ROB_ID_WIDTH - 1                  : 0]    o_exu_rob_rob_id_0,
    output  [31                                 : 0]    o_exu_rob_fence_src1,
    output  [31                                 : 0]    o_exu_rob_fence_src2,

    output                                              o_exu_rsv_wren_1,
    output  [`PRF_CODE_WIDTH - 1                : 0]    o_exu_rsv_wr_prf_code_1,
    output  [`PRF_DATA_WIDTH - 1                : 0]    o_exu_rsv_wr_dat_1,
    output                                              o_exu_rsv_busy_1,
    output                                              o_exu_rob_vld_1,
    output  [`ROB_ID_WIDTH - 1                  : 0]    o_exu_rob_rob_id_1,
    output  [`EXCEPTION_CODE_WIDTH - 1          : 0]    o_exu_rob_excp_code_1,
    output                                              o_exu_mis_flush,
    output  [`ROB_ID_WIDTH - 1                  : 0]    o_exu_mis_rob_id,
    output  [`CORE_PC_WIDTH - 1                 : 0]    o_exu_mis_addr,
    output                                              o_exu_iq_btac_vld,
    output                                              o_exu_iq_btac_taken,
    output                                              o_exu_iq_btac_new_br,
    output                                              o_exu_iq_type,
    output  [`CORE_PC_WIDTH - 1                 : 0]    o_exu_iq_btac_addr,
    output  [`CORE_PC_WIDTH - 1                 : 0]    o_exu_iq_btac_taddr,
    output  [1                                  : 0]    o_exu_iq_btac_idx,
    output  [`IQ_PHT_IDX_WIDTH - 1              : 0]    o_exu_iq_pht_idx,
    output  [1                                  : 0]    o_exu_iq_pht_status,
    output                                              o_exu_iq_len,
    output                                              o_exu_iq_tsucc, 

    output                                              o_exu_rsv_wren_2,
    output  [`PRF_CODE_WIDTH - 1                : 0]    o_exu_rsv_wr_prf_code_2,
    output  [`PRF_DATA_WIDTH - 1                : 0]    o_exu_rsv_wr_dat_2,
    output                                              o_exu_rsv_busy_2,
    output                                              o_exu_rob_vld_2,
    output  [`EXCEPTION_CODE_WIDTH - 1          : 0]    o_exu_rob_excp_code_2,
    output  [`ROB_ID_WIDTH - 1                  : 0]    o_exu_rob_rob_id_2,

    output                                              o_exu_rsv_wren_3,
    output  [`PRF_CODE_WIDTH - 1                : 0]    o_exu_rsv_wr_prf_code_3,
    output  [`PRF_DATA_WIDTH - 1                : 0]    o_exu_rsv_wr_dat_3,
    output                                              o_exu_rsv_busy_3,
    output                                              o_exu_rob_vld_3,
    output  [`EXCEPTION_CODE_WIDTH - 1          : 0]    o_exu_rob_excp_code_3,
    output  [`ROB_ID_WIDTH - 1                  : 0]    o_exu_rob_rob_id_3,
    output                                              o_exu_ls_flush,
    output  [`ROB_ID_WIDTH - 1                  : 0]    o_exu_ls_rob_id,
    output  [`CORE_PC_WIDTH - 1                 : 0]    o_exu_ls_addr,
    output                                              o_dtlb_mmu_vld,
    output  [`CORE_PC_WIDTH - 1                 : 0]    o_dtlb_mmu_vaddr,
    output                                              o_exu_mem_rd_vld,
    output  [`PHY_ADDR_WIDTH - 1                : 0]    o_exu_mem_rd_paddr,
    output                                              o_exu_mem_wr_vld,
    output  [`DCACHE_DATA_WIDTH - 1             : 0]    o_exu_mem_wdat,
    output  [`PHY_ADDR_WIDTH - 1                : 0]    o_exu_mem_wr_paddr,
    output                                              o_exu_dsp_s_ret,
    output                                              o_exu_rob_s_ret_done,

    input                                               clk,
    input                                               rst_n
);

//  ALU
alu_module alu ( 
    .i_csr_trap_flush     (i_csr_trap_flush),
    .i_exu_mis_flush      (o_exu_mis_flush),
    .i_exu_mis_rob_id     (o_exu_mis_rob_id),
    .i_exu_ls_flush       (o_exu_ls_flush),
    .i_exu_ls_rob_id      (o_exu_ls_rob_id),

    .i_rsv_exu_vld        (i_rsv_exu_vld_0),
    .i_rsv_exu_src1_vld   (i_rsv_exu_src1_vld_0),
    .i_rsv_exu_src1_dat   (i_rsv_exu_src1_dat_0),
    .i_rsv_exu_src2_vld   (i_rsv_exu_src2_vld_0),
    .i_rsv_exu_src2_dat   (i_rsv_exu_src2_dat_0),
    .i_rsv_exu_src3_vld   (i_rsv_exu_src3_vld_0),
    .i_rsv_exu_src3_dat   (i_rsv_exu_src3_dat_0),
    .i_rsv_exu_dst_vld    (i_rsv_exu_dst_vld_0),
    .i_rsv_exu_dst_code   (i_rsv_exu_dst_code_0),
    .i_rsv_exu_imm        (i_rsv_exu_imm_0),
    .i_rsv_exu_rob_id     (i_rsv_exu_rob_id_0),
    .i_rsv_exu_decinfo_bus(i_rsv_exu_decinfo_bus_0),
    .i_rsv_exu_len        (i_rsv_exu_len_0),
    .i_rob_exu_addr       (i_rob_exu_addr_0),
    .i_rsv_exu_excp_code  (i_rsv_exu_excp_code_0),
    .i_csr_exu_rdat       (i_csr_exu_rdat_0),
    .o_exu_csr_addr       (o_exu_csr_addr),
    .o_exu_csr_wren       (o_exu_csr_wren),
    .o_exu_csr_wdat       (o_exu_csr_wdat),
    .o_exu_rsv_wren       (o_exu_rsv_wren_0),
    .o_exu_rsv_wr_prf_code(o_exu_rsv_wr_prf_code_0),
    .o_exu_rsv_wdat       (o_exu_rsv_wr_dat_0),
    .o_exu_rsv_busy       (o_exu_rsv_busy_0),
    .o_exu_rob_vld        (o_exu_rob_vld_0),
    .o_exu_rob_excp_code  (o_exu_rob_excp_code_0),
    .o_exu_rob_done       (o_exu_rob_done_0),
    .o_exu_rob_rob_id     (o_exu_rob_rob_id_0),
    .o_exu_rob_fence_src1 (o_exu_rob_fence_src1),
    .o_exu_rob_fence_src2 (o_exu_rob_fence_src2),

    .clk                  (clk),
    .rst_n                (rst_n)
);

//  BJP
bjp_module bjp ( 
    .i_csr_trap_flush      (i_csr_trap_flush),
    .i_exu_ls_flush        (o_exu_ls_flush),
    .i_exu_ls_rob_id       (o_exu_ls_rob_id),

    .i_rsv_exu_vld         (i_rsv_exu_vld_1),
    .i_rsv_exu_src1_vld    (i_rsv_exu_src1_vld_1),
    .i_rsv_exu_src1_dat    (i_rsv_exu_src1_dat_1),
    .i_rsv_exu_src2_vld    (i_rsv_exu_src2_vld_1),
    .i_rsv_exu_src2_dat    (i_rsv_exu_src2_dat_1),
    .i_rsv_exu_src3_vld    (i_rsv_exu_src3_vld_1),
    .i_rsv_exu_src3_dat    (i_rsv_exu_src3_dat_1),
    .i_rsv_exu_imm         (i_rsv_exu_imm_1),
    .i_rsv_exu_decinfo_bus (i_rsv_exu_decinfo_bus_1),
    .i_rsv_exu_predinfo_bus(i_rsv_exu_predinfo_bus_1),
    .i_rsv_exu_len         (i_rsv_exu_len_1),
    .i_rsv_exu_rob_id      (i_rsv_exu_rob_id_1),
    .i_rsv_exu_excp_code   (i_rsv_exu_excp_code_1),
    .i_rob_exu_addr        (i_rob_exu_addr_1),
    .i_rob_exu_taddr       (i_rob_exu_taddr_1),

    .o_exu_rsv_wren        (o_exu_rsv_wren_1),
    .o_exu_rsv_wr_prf_code (o_exu_rsv_wr_prf_code_1),
    .o_exu_rsv_wr_dat      (o_exu_rsv_wr_dat_1),
    .o_exu_rob_vld         (o_exu_rob_vld_1),
    .o_exu_rob_rob_id      (o_exu_rob_rob_id_1),
    .o_exu_rob_excp_code   (o_exu_rob_excp_code_1),
    .o_exu_mis_flush       (o_exu_mis_flush),
    .o_exu_mis_rob_id      (o_exu_mis_rob_id),
    .o_exu_mis_addr        (o_exu_mis_addr),
    .o_exu_iq_btac_vld     (o_exu_iq_btac_vld),
    .o_exu_iq_btac_taken   (o_exu_iq_btac_taken),
    .o_exu_iq_btac_new_br  (o_exu_iq_btac_new_br),
    .o_exu_iq_type         (o_exu_iq_type),
    .o_exu_iq_btac_addr    (o_exu_iq_btac_addr),
    .o_exu_iq_btac_taddr   (o_exu_iq_btac_taddr),
    .o_exu_iq_btac_idx     (o_exu_iq_btac_idx),
    .o_exu_iq_pht_idx      (o_exu_iq_pht_idx),
    .o_exu_iq_pht_status   (o_exu_iq_pht_status),
    .o_exu_iq_len          (o_exu_iq_len),
    .o_exu_iq_tsucc        (o_exu_iq_tsucc),

    .clk                   (clk),
    .rst_n                 (rst_n)
);


//  MULDIV
exu_muldiv_module muldiv ( 
    .i_csr_trap_flush     (i_csr_trap_flush),
    .i_exu_mis_flush      (o_exu_mis_flush),
    .i_exu_mis_rob_id     (o_exu_mis_rob_id),
    .i_exu_ls_flush       (o_exu_ls_flush),
    .i_exu_ls_rob_id      (o_exu_ls_rob_id),

    .i_rsv_exu_vld        (i_rsv_exu_vld_2),
    .i_rsv_exu_src1_vld   (i_rsv_exu_src1_vld_2),
    .i_rsv_exu_src1_dat   (i_rsv_exu_src1_dat_2),
    .i_rsv_exu_src2_vld   (i_rsv_exu_src2_vld_2),
    .i_rsv_exu_src2_dat   (i_rsv_exu_src2_dat_2),
    .i_rsv_exu_src3_vld   (i_rsv_exu_src3_vld_2),
    .i_rsv_exu_src3_dat   (i_rsv_exu_src3_dat_2),
    .i_rsv_exu_dst_vld    (i_rsv_exu_dst_vld_2),
    .i_rsv_exu_dst_code   (i_rsv_exu_dst_code_2),
    .i_rsv_exu_decinfo_bus(i_rsv_exu_decinfo_bus_2),
    .i_rsv_exu_excp_code  (i_rsv_exu_excp_code_2),
    .i_rsv_exu_rob_id     (i_rsv_exu_rob_id_2),
    
    .o_exu_rsv_wren       (o_exu_rsv_wren_2),
    .o_exu_rsv_wr_prf_code(o_exu_rsv_wr_prf_code_2),
    .o_exu_rsv_wr_dat     (o_exu_rsv_wr_dat_2),
    .o_exu_rsv_busy       (o_exu_rsv_busy_2),
    .o_exu_rob_vld        (o_exu_rob_vld_2),
    .o_exu_rob_excp_code  (o_exu_rob_excp_code_2),
    .o_exu_rob_rob_id     (o_exu_rob_rob_id_2),

    .clk                  (clk),
    .rst_n                (rst_n)
);


//  AGU
exu_agu_module agu ( 
    .i_csr_trap_flush       (i_csr_trap_flush),
    .i_exu_mis_flush        (i_exu_mis_flush),
    .i_exu_mis_rob_id       (i_exu_mis_rob_id),
    .i_csr_rv_mode          (i_csr_rv_mode),
    .i_csr_mmu_satp         (i_csr_mmu_satp),

    .i_dsp_rsv_vld          (i_dsp_rsv_vld),
    .i_dsp_rsv_rob_id_0     (i_dsp_rsv_rob_id_0),
    .i_dsp_rsv_ld_vld_0     (i_dsp_rsv_ld_vld_0),
    .i_dsp_rsv_ld_id_0      (i_dsp_rsv_ld_id_0),
    .i_dsp_rsv_st_vld_0     (i_dsp_rsv_st_vld_0),
    .i_dsp_rsv_st_id_0      (i_dsp_rsv_st_id_0),
    .i_dsp_rsv_dst_vld_0    (i_dsp_rsv_dst_vld_0),
    .i_dsp_rsv_dst_code_0   (i_dsp_rsv_dst_code_0),
    .i_dsp_rsv_decinfo_bus_0(i_dsp_rsv_decinfo_bus_0),
    .i_dsp_rsv_rob_id_1     (i_dsp_rsv_rob_id_1),
    .i_dsp_rsv_ld_vld_1     (i_dsp_rsv_ld_vld_1),
    .i_dsp_rsv_ld_id_1      (i_dsp_rsv_ld_id_1),
    .i_dsp_rsv_st_vld_1     (i_dsp_rsv_st_vld_1),
    .i_dsp_rsv_st_id_1      (i_dsp_rsv_st_id_1),
    .i_dsp_rsv_dst_vld_1    (i_dsp_rsv_dst_vld_1),
    .i_dsp_rsv_dst_code_1   (i_dsp_rsv_dst_code_1),
    .i_dsp_rsv_decinfo_bus_1(i_dsp_rsv_decinfo_bus_1),
    .i_dsp_rsv_rob_id_2     (i_dsp_rsv_rob_id_2),
    .i_dsp_rsv_ld_vld_2     (i_dsp_rsv_ld_vld_2),
    .i_dsp_rsv_ld_id_2      (i_dsp_rsv_ld_id_2),
    .i_dsp_rsv_st_vld_2     (i_dsp_rsv_st_vld_2),
    .i_dsp_rsv_st_id_2      (i_dsp_rsv_st_id_2),
    .i_dsp_rsv_dst_vld_2    (i_dsp_rsv_dst_vld_2),
    .i_dsp_rsv_dst_code_2   (i_dsp_rsv_dst_code_2),
    .i_dsp_rsv_decinfo_bus_2(i_dsp_rsv_decinfo_bus_2),
    .i_dsp_rsv_rob_id_3     (i_dsp_rsv_rob_id_3),
    .i_dsp_rsv_ld_vld_3     (i_dsp_rsv_ld_vld_3),
    .i_dsp_rsv_ld_id_3      (i_dsp_rsv_ld_id_3),
    .i_dsp_rsv_st_vld_3     (i_dsp_rsv_st_vld_3),
    .i_dsp_rsv_st_id_3      (i_dsp_rsv_st_id_3),
    .i_dsp_rsv_dst_vld_3    (i_dsp_rsv_dst_vld_3),
    .i_dsp_rsv_dst_code_3   (i_dsp_rsv_dst_code_3),
    .i_dsp_rsv_decinfo_bus_3(i_dsp_rsv_decinfo_bus_3),
    .i_dsp_exu_ld_dsp_ptr   (i_dsp_exu_ld_dsp_ptr),
    .i_dsp_exu_ld_ret_ptr   (i_dsp_exu_ld_ret_ptr),
    .i_dsp_exu_st_dsp_ptr   (i_dsp_exu_st_dsp_ptr),
    .i_dsp_exu_st_ret_ptr   (i_dsp_exu_st_ret_ptr),
    .i_dsp_exu_st_ret_cptr  (i_dsp_exu_st_ret_cptr),

    .i_rob_exu_ret_vld      (i_rob_exu_ret_vld),
    .i_rob_exu_ret_ld_vld_0 (i_rob_exu_ret_ld_vld_0),
    .i_rob_exu_ret_ld_id_0  (i_rob_exu_ret_ld_id_0),
    .i_rob_exu_ret_st_vld_0 (i_rob_exu_ret_st_vld_0),
    .i_rob_exu_ret_st_id_0  (i_rob_exu_ret_st_id_0),
    .i_rob_exu_ret_ld_vld_1 (i_rob_exu_ret_ld_vld_1),
    .i_rob_exu_ret_ld_id_1  (i_rob_exu_ret_ld_id_1),
    .i_rob_exu_ret_st_vld_1 (i_rob_exu_ret_st_vld_1),
    .i_rob_exu_ret_st_id_1  (i_rob_exu_ret_st_id_1),
    .i_rob_exu_ret_ld_vld_2 (i_rob_exu_ret_ld_vld_2),
    .i_rob_exu_ret_ld_id_2  (i_rob_exu_ret_ld_id_2),
    .i_rob_exu_ret_st_vld_2 (i_rob_exu_ret_st_vld_2),
    .i_rob_exu_ret_st_id_2  (i_rob_exu_ret_st_id_2),
    .i_rob_exu_ret_ld_vld_3 (i_rob_exu_ret_ld_vld_3),
    .i_rob_exu_ret_ld_id_3  (i_rob_exu_ret_ld_id_3),
    .i_rob_exu_ret_st_vld_3 (i_rob_exu_ret_st_vld_3),
    .i_rob_exu_ret_st_id_3  (i_rob_exu_ret_st_id_3),
    .i_rob_exu_ls_addr      (i_rob_exu_ls_addr),
    .i_rob_dtlb_flush       (i_rob_dtlb_flush),
    .i_rob_dtlb_src1        (i_rob_dtlb_src1),
    .i_rob_dtlb_src2        (i_rob_dtlb_src2),

    .i_rsv_exu_vld          (i_rsv_exu_vld),
    .i_rsv_exu_src1_vld     (i_rsv_exu_src1_vld_3),
    .i_rsv_exu_src1_dat     (i_rsv_exu_src1_dat_3),
    .i_rsv_exu_src2_vld     (i_rsv_exu_src2_vld_3),
    .i_rsv_exu_src2_dat     (i_rsv_exu_src2_dat_3),
    .i_rsv_exu_src3_vld     (i_rsv_exu_src3_vld_3),
    .i_rsv_exu_src3_dat     (i_rsv_exu_src3_dat_3),
    .i_rsv_exu_dst_vld      (i_rsv_exu_dst_vld_3),
    .i_rsv_exu_dst_code     (i_rsv_exu_dst_code_3),
    .i_rsv_exu_rob_id       (i_rsv_exu_rob_id_3),
    .i_rsv_exu_ld_vld       (i_rsv_exu_ld_vld_3),
    .i_rsv_exu_ld_id        (i_rsv_exu_ld_id_3),
    .i_rsv_exu_st_vld       (i_rsv_exu_st_vld_3),
    .i_rsv_exu_st_id        (i_rsv_exu_st_id_3),
    .i_rsv_exu_decinfo_bus  (i_rsv_exu_decinfo_bus_3),
    .i_rsv_exu_imm          (i_rsv_exu_imm_3),

    .i_mmu_busy             (i_mmu_busy),
    .i_mmu_dtlb_vld         (i_mmu_dtlb_vld),
    .i_mmu_dtlb_tlb         (i_mmu_dtlb_tlb),
    .i_mmu_dtlb_excp_code   (i_mmu_dtlb_excp_code),
    .i_mmu_dcache_vld       (i_mmu_dcache_vld),
    .i_mmu_dcache_dat       (i_mmu_dcache_dat),
    .i_mmu_exu_done         (i_mmu_exu_done),

    .o_exu_rsv_wren         (o_exu_rsv_wren_3),
    .o_exu_rsv_wr_prf_code  (o_exu_rsv_wr_prf_code_3),
    .o_exu_rsv_wr_dat       (o_exu_rsv_wr_dat_3),
    .o_exu_rsv_busy         (o_exu_rsv_busy_3),
    .o_exu_rob_vld          (o_exu_rob_vld_3),
    .o_exu_rob_excp_code    (o_exu_rob_excp_code_3),
    .o_exu_rob_rob_id       (o_exu_rob_rob_id_3),
    .o_exu_ls_flush         (o_exu_ls_flush),
    .o_exu_ls_rob_id        (o_exu_ls_rob_id),
    .o_exu_ls_addr          (o_exu_ls_addr),
    .o_dtlb_mmu_vld         (o_dtlb_mmu_vld),
    .o_dtlb_mmu_vaddr       (o_dtlb_mmu_vaddr),
    .o_exu_mem_rd_vld       (o_exu_mem_rd_vld),
    .o_exu_mem_rd_paddr     (o_exu_mem_rd_paddr),
    .o_exu_mem_wr_vld       (o_exu_mem_wr_vld),
    .o_exu_mem_wdat         (o_exu_mem_wdat),
    .o_exu_mem_wr_paddr     (o_exu_mem_wr_paddr),
    .o_exu_dsp_s_ret        (o_exu_dsp_s_ret),
    .o_exu_dsp_s_ret_done   (o_exu_dsp_s_ret_done),

    .clk                    (clk),
    .rst_n                  (rst_n)
);

endmodule   //  exu_top_module

`endif  /*  !__EXU_EXU_TOP_V__! */