`ifdef __EXU_EXU_DCACHE_V__

module exu_dcache_module (

);


endmodule   //  exu_dcache_module

`endif  /*  !__EXU_EXU_DCACHE_V__!  */